/*
This file creates the test bench for the systolic array method

The goal is to store a matrix in a bram in the Tb and then during the test itself call the systolic array method and see 
it work

The question is how to parametize the function!

*/